// Register File - Per-lane register file
// TODO: Implement per-lane register file
// - 32 registers × 32 bits (configurable)
// - Dual-port for read/write in same cycle
// - Register 0 hardwired to zero

module register_file (
    // TODO: Add module ports (clock, read_addr1, read_addr2, write_addr, write_data, read_data1, read_data2, write_en)
);

    // TODO: Implement register array
    // TODO: Implement dual-port read
    // TODO: Implement write port
    // TODO: Hardwire register 0 to zero

endmodule

