// RoCC Interface - Standard RoCC command decoder (core-agnostic)
// TODO: Implement RoCC interface following standard RoCC spec
// - io.cmd.* (command interface)
// - io.resp.* (response interface)
// - io.mem.* (memory interface)
// - Custom instructions: kernel_start, set_mask, get_status

module rocc_interface (
    // TODO: Add RoCC interface ports
);

    // TODO: Implement command decoding
    // TODO: Implement kernel descriptor handling
    // TODO: Implement memory request handling
    // TODO: Implement status reporting

endmodule

