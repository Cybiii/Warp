// Warp Controller Testbench
// TODO: Implement warp controller testbench
// - Test FSM transitions (IDLE, LOAD, EXECUTE, STALL, DONE)
// - Test control flow
// - Test stall conditions

`timescale 1ns/1ps

module tb_warp_controller;

    // TODO: Add testbench signals
    // TODO: Instantiate warp_controller
    // TODO: Test FSM state transitions
    // TODO: Test control signals

    initial begin
        // TODO: Test IDLE -> LOAD transition
        // TODO: Test LOAD -> EXECUTE transition
        // TODO: Test EXECUTE -> STALL transition
        // TODO: Test STALL -> EXECUTE transition
        // TODO: Test EXECUTE -> DONE transition
        $finish;
    end

endmodule

